library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
entity DigitalClock is port(
	soundclk:in std_logic;	--����ʱ��Ƶ�� ĿǰΪ100K
	turnOn:in std_logic;		--�����ź� ����Ч��Ĭ��Ӧ��Ϊ0 
	spk:out std_logic			--������Ƶ�����
);
end entity;

architecture behav of DigitalClock is
signal clk: std_logic_vector(15 downto 0):="0000000000000000";		--��Ƶ���ʱ�������
signal reset: std_logic:='0'; 	--��λ�ź� ����Ч
signal waveout: std_logic;       --����ź�
signal freq: std_logic_vector(7 downto 0);
signal soundcnt:std_logic_vector(7 downto 0);				--clk���ڼ����� 
signal dotcnt:std_logic_vector(3 downto 0) ;		--������ż���
signal songcnt:std_logic_vector(2 downto 0);  	--����ѭ����������

constant spkout:std_logic_vector(15 downto 0):="1001110001000000"; --������10Hz,10K
constant do:std_logic_vector(7 downto 0):="10111111";	--do��Ƶ��100KHz/261.6Hz/2=191.1(��������)��������10111111
constant re:std_logic_vector(7 downto 0):="10101010";	--re��Ƶ��293.7Hz������ͬ��
constant mi:std_logic_vector(7 downto 0):="10010111";	--mi��Ƶ��329.6Hz������ͬ��
constant fa:std_logic_vector(7 downto 0):="10001111";	--fa��Ƶ��349.2Hz������ͬ��
constant so:std_logic_vector(7 downto 0):="01111111";	--so��Ƶ��392Hz������ͬ��
constant la:std_logic_vector(7 downto 0):="01110001";	--la��Ƶ��440Hz������ͬ��
constant si:std_logic_vector(7 downto 0):="01100101";	--la��Ƶ��493.9Hz������ͬ��
constant non:std_logic_vector(7 downto 0):="00000000"; --��Ƶ��ֵ

begin
	spk <= waveout;

	process(soundclk,turnOn)
	begin
		if (soundclk'event and soundclk='1') then
		
		--��������
			if turnOn = '1' then reset <= '1'; songcnt <= "000"; dotcnt <= "0000";		--��ʼ����
			end if;
				--���ӵ�����(��ǰ)
			if clk = spkout 		--����������ﵽ���ڣ���ʼ��������
				then clk <= "0000000000000000";
			
				if songcnt = "100" then freq <= non; songcnt <= "000"; reset <= '0';		--����ѭ�������Ѵֹͣ
				end if;
			
				if reset = '1' then																		--������ڲ���״̬����ʼ��������
					case dotcnt is			
						when "0000" => freq <= do; dotcnt <= dotcnt + 1;
						when "0001" => freq <= re; dotcnt <= dotcnt + 1;
						when "0010" => freq <= mi; dotcnt <= dotcnt + 1;
						when "0011" => freq <= do; dotcnt <= dotcnt + 1;
						when "0100" => freq <= do; dotcnt <= dotcnt + 1;
						when "0101" => freq <= re; dotcnt <= dotcnt + 1;
						when "0110" => freq <= mi; dotcnt <= dotcnt + 1;
						when "0111" => freq <= do; dotcnt <= dotcnt + 1;
						when "1000" => freq <= mi; dotcnt <= dotcnt + 1;
						when "1001" => freq <= fa; dotcnt <= dotcnt + 1;
						when "1010" => freq <= so; dotcnt <= dotcnt + 1;
						when "1011" => freq <= non; dotcnt <= dotcnt + 1;
						when "1100" => freq <= mi; dotcnt <= dotcnt + 1;
						when "1101" => freq <= fa; dotcnt <= dotcnt + 1;
						when "1110" => freq <= so;dotcnt <= "0000"; songcnt <= songcnt + 1;
						when others => freq <= fa; dotcnt <= "0000"; songcnt <= songcnt + 1;
					end case;
				end if;
			else clk <= clk + 1;
			end if;
		--����
		
		--��Ƶ���
			if reset = '1' then 
				if freq = non 			--û����������
					then waveout <= '0';			--��������������������
				else
					if soundcnt = freq 		--�������ﵽ����
						then soundcnt <= "00000000";
						waveout <= not waveout;	--���ȡ�����������
					else soundcnt <= soundcnt + 1;
					end if;
				end if;
			
			else --��λ�ź���Чʱ
				waveout <= '0';
				soundcnt <= "00000000";
			end if;
		--����
		end if;
	end process;
end architecture;